magic
tech sky130A
magscale 1 2
timestamp 1622200441
<< metal1 >>
rect 150 2602 350 2792
rect -58 2598 566 2602
rect -58 2134 570 2598
rect -266 2032 286 2074
rect -264 1754 -230 2032
rect 492 2002 570 2134
rect 90 1962 570 2002
rect 182 1792 630 1838
rect -264 1732 388 1754
rect -262 1696 388 1732
rect -790 1438 -590 1510
rect -262 1438 -204 1696
rect -790 1380 -204 1438
rect -790 1310 -590 1380
rect -262 1147 -204 1380
rect 580 1445 630 1792
rect 1128 1445 1328 1524
rect 580 1395 1328 1445
rect -262 1089 291 1147
rect -262 718 -204 1089
rect 580 1054 630 1395
rect 1128 1324 1328 1395
rect 184 1006 630 1054
rect 176 796 570 798
rect 86 760 570 796
rect 176 756 570 760
rect -262 689 383 718
rect -258 667 383 689
rect 478 630 566 756
rect -60 282 566 630
rect -60 274 518 282
rect 180 88 380 274
use sky130_fd_pr__nfet_01v8_N39HBR  XM1
timestamp 1622193717
transform 1 0 258 0 1 907
box -311 -360 311 360
use sky130_fd_pr__pfet_01v8_KG2LE3  XM2
timestamp 1622193717
transform 1 0 257 0 1 1889
box -311 -319 311 319
<< labels >>
flabel metal1 -790 1310 -590 1510 0 FreeSans 256 0 0 0 in
port 1 nsew
flabel metal1 1128 1324 1328 1524 0 FreeSans 256 0 0 0 out
port 0 nsew
flabel metal1 180 88 380 288 0 FreeSans 256 0 0 0 vss
port 2 nsew
flabel metal1 150 2592 350 2792 0 FreeSans 256 0 0 0 vdd
port 3 nsew
<< end >>
